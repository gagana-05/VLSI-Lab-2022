* nmos characteristics varying width

* include model files
.include ./t14y_tsmc_025_level3.txt

*netlist
*model instance 
m1 Vdd in Vss 0 cmosn w=0.5u l=1u

* voltage inputs
v_dd Vdd 0 3.3
v_ss Vss 0 0
v_in in 0 3.3

* plotting outputs for various widths
.control 
dc v_in 0 3.3 1 v_dd 0 3.3 1
foreach len 0.5u 10u
 alter m1 l=$len
run 
end
.endc

.control
foreach iter 1 2 
setplot dc$iter
plot -v_dd#branch
end
.endc
.end