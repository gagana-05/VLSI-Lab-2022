magic
tech scmos
timestamp 1668001487
<< nwell >>
rect 0 43 49 74
<< polysilicon >>
rect 7 63 9 65
rect 24 63 26 65
rect 41 63 43 65
rect 7 25 9 43
rect 24 25 26 43
rect 41 25 43 43
rect 7 11 9 13
rect 24 11 26 13
rect 41 11 43 13
<< ndiffusion >>
rect 1 22 7 25
rect 1 18 2 22
rect 6 18 7 22
rect 1 13 7 18
rect 9 22 24 25
rect 9 18 10 22
rect 14 18 24 22
rect 9 13 24 18
rect 26 22 41 25
rect 26 18 27 22
rect 31 18 41 22
rect 26 13 41 18
rect 43 22 49 25
rect 43 18 44 22
rect 48 18 49 22
rect 43 13 49 18
<< pdiffusion >>
rect 1 59 7 63
rect 1 55 2 59
rect 6 55 7 59
rect 1 43 7 55
rect 9 59 15 63
rect 9 55 10 59
rect 14 55 15 59
rect 9 43 15 55
rect 18 59 24 63
rect 18 55 19 59
rect 23 55 24 59
rect 18 43 24 55
rect 26 59 32 63
rect 26 55 27 59
rect 31 55 32 59
rect 26 43 32 55
rect 35 59 41 63
rect 35 55 36 59
rect 40 55 41 59
rect 35 43 41 55
rect 43 59 49 63
rect 43 55 44 59
rect 48 55 49 59
rect 43 43 49 55
<< metal1 >>
rect 1 73 49 74
rect 1 69 2 73
rect 6 69 49 73
rect 1 66 49 69
rect 2 59 6 66
rect 14 55 19 59
rect 31 55 36 59
rect 44 32 48 55
rect 10 28 48 32
rect 10 22 14 28
rect 2 10 6 18
rect 27 10 31 18
rect 44 10 48 18
rect 2 6 49 10
rect 6 2 27 6
rect 31 2 44 6
rect 48 2 49 6
rect 2 0 49 2
<< ntransistor >>
rect 7 13 9 25
rect 24 13 26 25
rect 41 13 43 25
<< ptransistor >>
rect 7 43 9 63
rect 24 43 26 63
rect 41 43 43 63
<< polycontact >>
rect 3 35 7 39
rect 20 35 24 39
rect 37 35 41 39
<< ndcontact >>
rect 2 18 6 22
rect 10 18 14 22
rect 27 18 31 22
rect 44 18 48 22
<< pdcontact >>
rect 2 55 6 59
rect 10 55 14 59
rect 19 55 23 59
rect 27 55 31 59
rect 36 55 40 59
rect 44 55 48 59
<< psubstratepcontact >>
rect 2 2 6 6
rect 27 2 31 6
rect 44 2 48 6
<< nsubstratencontact >>
rect 2 69 6 73
<< labels >>
rlabel psubstratepcontact 30 5 30 5 1 Vss
rlabel metal1 26 70 26 70 5 Vdd
rlabel polycontact 22 36 22 36 1 b
rlabel metal1 46 37 46 37 7 out
rlabel polycontact 39 37 39 37 1 c
rlabel polycontact 4 37 4 37 3 a
<< end >>
