* nmos characteristics

* include model files
.include ./t14y_tsmc_025_level1.txt

*netlist
* model instance 
m1 Vdd in Vss Vsb RITSUBN1 w=0.5u l=1u 

* voltage inputs
v_dd Vdd 0 3.3
v_ss Vss 0 0
v_sb Vsb 0 0

v_in in 0 3.3

.control 
* dc v_in 0 3.3 0.1 v_dd 0 3.3 1
dc v_dd 0 3.3 0.1 v_sb 0 3.3 1
run 
setplot dc1
plot -v_dd#branch

* dc v_dd 0 3.3 0.1 v_in 0 3.3 1
dc v_in 0 3.3 0.1 v_sb 0 3.3 1
run 
setplot dc2
plot -v_dd#branch
.endc

* .control
* foreach tem 10 25 50
* 	alter m1 TEMP=$tem	
* 	dc v_in 0 3.3 0.1 v_dd 0 3.3 1
*     run	
* end
* * alter m1 TEMP=27
* .endc

* .control
* foreach l 1 10 50
* 	altermod m1 LAMBDA=$l
* 	dc v_dd 0 3.3 0.1 v_in 0 3.3 1
* 	run
* end
* alter m1 LAMBDA= 0.031
* .endc
* .control
* foreach iter 1 2 3
* setplot dc$iter
* plot -v_dd#branch
* end
* .endc



.end