magic
tech scmos
timestamp 1667987679
<< nwell >>
rect 0 44 79 75
rect 39 43 79 44
<< polysilicon >>
rect 7 64 9 66
rect 24 64 26 66
rect 58 64 60 66
rect 7 26 9 44
rect 24 26 26 44
rect 58 32 60 44
rect 7 12 9 14
rect 24 12 26 14
rect 58 12 60 14
<< ndiffusion >>
rect 1 23 7 26
rect 1 19 2 23
rect 6 19 7 23
rect 1 14 7 19
rect 9 23 24 26
rect 9 19 10 23
rect 14 19 24 23
rect 9 14 24 19
rect 26 23 32 26
rect 26 19 27 23
rect 31 19 32 23
rect 26 14 32 19
rect 52 24 58 32
rect 52 20 53 24
rect 57 20 58 24
rect 52 14 58 20
rect 60 24 66 32
rect 60 20 61 24
rect 65 20 66 24
rect 60 14 66 20
<< pdiffusion >>
rect 1 60 7 64
rect 1 56 2 60
rect 6 56 7 60
rect 1 44 7 56
rect 9 60 15 64
rect 9 56 10 60
rect 14 56 15 60
rect 9 44 15 56
rect 18 60 24 64
rect 18 56 19 60
rect 23 56 24 60
rect 18 44 24 56
rect 26 60 32 64
rect 26 56 27 60
rect 31 56 32 60
rect 26 44 32 56
rect 52 59 58 64
rect 52 55 53 59
rect 57 55 58 59
rect 52 44 58 55
rect 60 59 66 64
rect 60 55 61 59
rect 65 55 66 59
rect 60 44 66 55
<< metal1 >>
rect 1 74 76 75
rect 1 70 2 74
rect 6 72 76 74
rect 6 70 53 72
rect 1 68 53 70
rect 57 68 76 72
rect 1 67 76 68
rect 2 60 6 67
rect 14 56 19 60
rect 31 56 37 60
rect 33 39 37 56
rect 53 59 57 67
rect 33 35 54 39
rect 33 33 37 35
rect 10 30 37 33
rect 10 23 14 30
rect 61 24 65 55
rect 2 11 6 19
rect 27 11 31 19
rect 53 11 57 20
rect 2 9 77 11
rect 2 7 53 9
rect 6 3 19 7
rect 23 5 53 7
rect 57 5 77 9
rect 23 3 77 5
rect 2 1 77 3
<< ntransistor >>
rect 7 14 9 26
rect 24 14 26 26
rect 58 14 60 32
<< ptransistor >>
rect 7 44 9 64
rect 24 44 26 64
rect 58 44 60 64
<< polycontact >>
rect 3 32 7 36
rect 20 36 24 40
rect 54 35 58 39
<< ndcontact >>
rect 2 19 6 23
rect 10 19 14 23
rect 27 19 31 23
rect 53 20 57 24
rect 61 20 65 24
<< pdcontact >>
rect 2 56 6 60
rect 10 56 14 60
rect 19 56 23 60
rect 27 56 31 60
rect 53 55 57 59
rect 61 55 65 59
<< psubstratepcontact >>
rect 2 3 6 7
rect 19 3 23 7
rect 53 5 57 9
<< nsubstratencontact >>
rect 2 70 6 74
rect 53 68 57 72
<< labels >>
rlabel metal1 63 37 63 37 1 out
rlabel metal1 69 71 69 71 5 Vdd
rlabel metal1 70 6 70 6 1 Vss
rlabel polycontact 4 34 4 34 3 a
rlabel polycontact 22 37 22 37 1 b
<< end >>
