* SPICE3 file created from or.ext - technology: scmos

.option scale=1u
.include ./t14y_tsmc_025_level3.txt

M1000 out a_9_14# Vdd Vdd cmosp w=20 l=2
+  ad=120 pd=52 as=240 ps=104
M1001 a_9_14# b a_9_44# Vdd cmosp w=20 l=2
+  ad=120 pd=52 as=240 ps=104
M1002 out a_9_14# Vss 0 cmosn w=18 l=2
+  ad=108 pd=48 as=252 ps=120
M1003 Vss b a_9_14# 0 cmosn w=12 l=2
+  ad=0 pd=0 as=180 ps=54
M1004 a_9_44# a Vdd Vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 a_9_14# a Vss 0 cmosn w=12 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_9_14# Vdd 4.39fF
C1 Vss 0 34.69fF
C2 out 0 2.07fF
C3 a_9_14# 0 14.38fF
C4 b 0 6.50fF
C5 a 0 6.50fF

* voltage input
v_dd Vdd 0 3.3
v_ss Vss 0 0 

v_ina a 0 pulse(0 3.3 0 0.1n 0 50n 100n)
v_inb b 0 pulse(0 3.3 0 0.1n 0 100n 200n)

* output
.control
tran 0.1n 200n
setplot tran1
plot b a
plot out
plot b a out
.endc
.end
