* SPICE3 file created from nand.ext - technology: scmos

.option scale=1u
.include ./t14y_tsmc_025_level3.txt

M1000 Vdd c out Vdd cmosp w=7 l=2
+  ad=126 pd=78 as=126 ps=78
M1001 a_8_18# a Vss Gnd cmosn w=7 l=2
+  ad=84 pd=52 as=42 ps=26
M1002 out b Vdd Vdd cmosp w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 out a Vdd Vdd cmosp w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 out c a_25_18# Gnd cmosn w=7 l=2
+  ad=42 pd=26 as=77 ps=50
M1005 a_25_18# b a_8_18# Gnd cmosn w=7 l=2
+  ad=0 pd=0 as=0 ps=0
C0 Vss Gnd 21.90fF
C1 out Gnd 10.43fF
C2 c Gnd 7.22fF
C3 b Gnd 7.22fF
C4 a Gnd 7.22fF

* voltage input
v_dd Vdd 0 3.3
v_ss Vss 0 0 

v_ina a 0 3.3 pulse(0 3.3 0 0.1n 0 20n 40n)
v_inb b 0 3.3 pulse(0 3.3 0 0.1n 0 40n 80n)
v_inc c 0 3.3 pulse(0 3.3 0 0.1n 0 80n 160n)

* output
.control
tran 1n 200n
setplot tran1
plot c b a
plot out
.endc
.end
