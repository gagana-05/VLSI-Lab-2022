magic
tech scmos
timestamp 1668151013
<< nwell >>
rect -4 46 48 66
<< polysilicon >>
rect 6 53 8 55
rect 23 53 25 55
rect 40 53 42 55
rect 6 25 8 46
rect 23 25 25 46
rect 40 25 42 46
rect 6 16 8 18
rect 23 16 25 18
rect 40 16 42 18
<< ndiffusion >>
rect 0 24 6 25
rect 0 20 1 24
rect 5 20 6 24
rect 0 18 6 20
rect 8 24 14 25
rect 8 20 9 24
rect 13 20 14 24
rect 8 18 14 20
rect 17 24 23 25
rect 17 20 18 24
rect 22 20 23 24
rect 17 18 23 20
rect 25 24 30 25
rect 25 20 26 24
rect 25 18 30 20
rect 34 24 40 25
rect 34 20 35 24
rect 39 20 40 24
rect 34 18 40 20
rect 42 24 48 25
rect 42 20 43 24
rect 47 20 48 24
rect 42 18 48 20
<< pdiffusion >>
rect 0 51 6 53
rect 0 47 1 51
rect 5 47 6 51
rect 0 46 6 47
rect 8 51 14 53
rect 8 47 9 51
rect 13 47 14 51
rect 8 46 14 47
rect 17 51 23 53
rect 17 47 18 51
rect 22 47 23 51
rect 17 46 23 47
rect 25 51 31 53
rect 25 47 26 51
rect 30 47 31 51
rect 25 46 31 47
rect 34 51 40 53
rect 34 47 35 51
rect 39 47 40 51
rect 34 46 40 47
rect 42 51 48 53
rect 42 47 43 51
rect 47 47 48 51
rect 42 46 48 47
<< metal1 >>
rect 0 63 48 64
rect 0 59 1 63
rect 5 59 18 63
rect 22 59 43 63
rect 47 59 48 63
rect 0 56 48 59
rect 1 51 5 56
rect 18 51 22 56
rect 43 51 47 56
rect 9 40 13 47
rect 26 40 30 47
rect 35 40 39 47
rect 9 36 47 40
rect 43 24 47 36
rect 13 20 18 24
rect 30 20 35 24
rect 1 15 5 20
rect 1 12 48 15
rect 5 8 48 12
rect 1 5 48 8
<< ntransistor >>
rect 6 18 8 25
rect 23 18 25 25
rect 40 18 42 25
<< ptransistor >>
rect 6 46 8 53
rect 23 46 25 53
rect 40 46 42 53
<< polycontact >>
rect 2 33 6 37
rect 19 29 23 33
rect 36 29 40 33
<< ndcontact >>
rect 1 20 5 24
rect 9 20 13 24
rect 18 20 22 24
rect 26 20 30 24
rect 35 20 39 24
rect 43 20 47 24
<< pdcontact >>
rect 1 47 5 51
rect 9 47 13 51
rect 18 47 22 51
rect 26 47 30 51
rect 35 47 39 51
rect 43 47 47 51
<< psubstratepcontact >>
rect 1 8 5 12
<< nsubstratencontact >>
rect 1 59 5 63
rect 18 59 22 63
rect 43 59 47 63
<< labels >>
rlabel polycontact 22 31 22 31 1 b
rlabel polycontact 4 35 4 35 3 a
rlabel metal1 45 31 45 31 7 out
rlabel polycontact 38 31 38 31 1 c
rlabel metal1 14 61 14 61 5 Vdd
rlabel metal1 14 10 14 10 1 Vss
<< end >>
