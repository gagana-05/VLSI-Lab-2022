* nmos characteristics varying length

* include model files
.include ./t14y_tsmc_025_level3.txt

*netlist
*model instance 
m1 Vdd in Vss 0 cmosn w=0.5u l=1u

* voltage inputs
v_dd Vdd 0 3.3
v_ss Vss 0 0
v_in in 0 3.3

* plotting outputs for various lengths
.control 
foreach len 0.5u 1u 2u 10u
 alter m1 l=$len
 dc v_dd 0 3.3 0.1 v_in 0 3.3 1
run 
end
.endc

.control
foreach iter 1 2 3 4
setplot dc$iter
plot -v_dd#branch
end
.endc
.end