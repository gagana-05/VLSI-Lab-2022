magic
tech scmos
timestamp 1667983989
<< polysilicon >>
rect 6 -3 8 -1
rect 6 -35 8 -23
rect 6 -55 8 -53
<< ndiffusion >>
rect 0 -43 6 -35
rect 0 -47 1 -43
rect 5 -47 6 -43
rect 0 -53 6 -47
rect 8 -43 14 -35
rect 8 -47 9 -43
rect 13 -47 14 -43
rect 8 -53 14 -47
<< pdiffusion >>
rect 0 -8 6 -3
rect 0 -12 1 -8
rect 5 -12 6 -8
rect 0 -23 6 -12
rect 8 -8 14 -3
rect 8 -12 9 -8
rect 13 -12 14 -8
rect 8 -23 14 -12
<< metal1 >>
rect 0 5 24 8
rect 0 1 1 5
rect 5 1 24 5
rect 0 0 24 1
rect 1 -8 5 0
rect 9 -43 13 -12
rect 1 -56 5 -47
rect 0 -58 25 -56
rect 0 -62 1 -58
rect 5 -62 25 -58
rect 0 -66 25 -62
<< ntransistor >>
rect 6 -53 8 -35
<< ptransistor >>
rect 6 -23 8 -3
<< polycontact >>
rect 2 -32 6 -28
<< ndcontact >>
rect 1 -47 5 -43
rect 9 -47 13 -43
<< pdcontact >>
rect 1 -12 5 -8
rect 9 -12 13 -8
<< psubstratepcontact >>
rect 1 -62 5 -58
<< nsubstratencontact >>
rect 1 1 5 5
<< labels >>
rlabel metal1 11 -30 11 -30 1 out
rlabel polycontact 4 -30 4 -30 3 a
rlabel metal1 17 4 17 4 5 Vdd
rlabel metal1 18 -61 18 -61 1 Vss
<< end >>
