* SPICE3 file created from gagana_joshua.ext - technology: scmos

.option scale=1u

M1000 out in Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1001 out in Vss Gnd nfet w=10 l=2
+  ad=50 pd=30 as=50 ps=30
C0 Vss Gnd 4.98fF
C1 out Gnd 2.07fF
C2 in Gnd 5.47fF
