magic
tech scmos
timestamp 1668018142
<< nwell >>
rect -4 42 48 76
<< polysilicon >>
rect 6 63 8 65
rect 23 63 25 65
rect 40 63 42 65
rect 6 25 8 43
rect 23 25 25 43
rect 40 25 42 43
rect 6 11 8 13
rect 23 11 25 13
rect 40 11 42 13
<< ndiffusion >>
rect 0 24 6 25
rect 0 20 1 24
rect 5 20 6 24
rect 0 13 6 20
rect 8 24 14 25
rect 8 20 9 24
rect 13 20 14 24
rect 8 13 14 20
rect 17 24 23 25
rect 17 20 18 24
rect 22 20 23 24
rect 17 13 23 20
rect 25 24 30 25
rect 25 20 26 24
rect 25 13 30 20
rect 34 24 40 25
rect 34 20 35 24
rect 39 20 40 24
rect 34 13 40 20
rect 42 24 48 25
rect 42 20 43 24
rect 47 20 48 24
rect 42 13 48 20
<< pdiffusion >>
rect 0 61 6 63
rect 0 57 1 61
rect 5 57 6 61
rect 0 43 6 57
rect 8 61 23 63
rect 8 57 9 61
rect 13 57 18 61
rect 22 57 23 61
rect 8 43 23 57
rect 25 61 40 63
rect 25 57 33 61
rect 37 57 40 61
rect 25 43 40 57
rect 42 61 48 63
rect 42 57 43 61
rect 47 57 48 61
rect 42 43 48 57
<< metal1 >>
rect 0 73 48 74
rect 0 69 1 73
rect 5 69 18 73
rect 22 69 43 73
rect 47 69 48 73
rect 0 66 48 69
rect 1 61 5 66
rect 18 61 22 66
rect 43 61 47 66
rect 9 40 13 57
rect 33 40 37 57
rect 9 36 47 40
rect 43 24 47 36
rect 13 20 18 24
rect 30 20 35 24
rect 1 10 5 20
rect 1 7 48 10
rect 5 3 48 7
rect 1 0 48 3
<< ntransistor >>
rect 6 13 8 25
rect 23 13 25 25
rect 40 13 42 25
<< ptransistor >>
rect 6 43 8 63
rect 23 43 25 63
rect 40 43 42 63
<< polycontact >>
rect 2 33 6 37
rect 19 29 23 33
rect 36 29 40 33
<< ndcontact >>
rect 1 20 5 24
rect 9 20 13 24
rect 18 20 22 24
rect 26 20 30 24
rect 35 20 39 24
rect 43 20 47 24
<< pdcontact >>
rect 1 57 5 61
rect 9 57 13 61
rect 18 57 22 61
rect 33 57 37 61
rect 43 57 47 61
<< psubstratepcontact >>
rect 1 3 5 7
<< nsubstratencontact >>
rect 1 69 5 73
rect 18 69 22 73
rect 43 69 47 73
<< labels >>
rlabel polycontact 22 31 22 31 1 b
rlabel polycontact 4 35 4 35 3 a
rlabel metal1 14 71 14 71 5 Vdd
rlabel metal1 14 5 14 5 1 Vss
rlabel metal1 45 31 45 31 7 out
rlabel polycontact 38 31 38 31 1 c
<< end >>
