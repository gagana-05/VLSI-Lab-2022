* include the model files
*.include ./t14y_tsmc_025_level3.txt
  
* netlist
* m_instance_name drain_node gate_node source_node bulk_substrate_node model_name L=length W=width
m0 out in vss 0 nfet l=2u w=10u 
m1 out in vdd 0 pfet l=2u w=20u

* power sources excitation etc.
* v_instance_name posive_node negetive_node value
* supply voltages
Vgnd vss 0 dc 0
*Vdd vdd 0 dc 3.3

v_dd vdd 0 3.3
* input voltage source:
Vin in 0 dc 2.5 pulse(0 5 1n 0.1n 0.1n 2n 4n) 
tran 0.1n 200n
plot -v_dd#branch


.end
