* SPICE3 file created from or.ext - technology: scmos

.option scale=1u

M1000 out a_9_14# Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=240 ps=104
M1001 a_9_14# b a_9_44# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=240 ps=104
M1002 out a_9_14# Vss Gnd nfet w=18 l=2
+  ad=108 pd=48 as=252 ps=120
M1003 Vss b a_9_14# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=180 ps=54
M1004 a_9_44# a Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 a_9_14# a Vss Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_9_14# Vdd 4.39fF
C1 Vss Gnd 34.69fF
C2 out Gnd 2.07fF
C3 a_9_14# Gnd 14.38fF
C4 b Gnd 6.50fF
C5 a Gnd 6.50fF
