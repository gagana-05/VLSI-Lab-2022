magic
tech scmos
timestamp 1667986998
<< nwell >>
rect 1 -19 75 16
<< polysilicon >>
rect 10 2 12 4
rect 27 2 29 4
rect 52 2 54 4
rect 10 -36 12 -18
rect 27 -36 29 -18
rect 52 -30 54 -18
rect 10 -50 12 -48
rect 27 -50 29 -48
rect 52 -50 54 -48
<< ndiffusion >>
rect 4 -37 10 -36
rect 4 -41 5 -37
rect 9 -41 10 -37
rect 4 -48 10 -41
rect 12 -37 18 -36
rect 12 -41 13 -37
rect 17 -41 18 -37
rect 12 -48 18 -41
rect 21 -37 27 -36
rect 21 -41 22 -37
rect 26 -41 27 -37
rect 21 -48 27 -41
rect 29 -37 34 -36
rect 29 -41 30 -37
rect 29 -48 34 -41
rect 46 -38 52 -30
rect 46 -42 47 -38
rect 51 -42 52 -38
rect 46 -48 52 -42
rect 54 -38 60 -30
rect 54 -42 55 -38
rect 59 -42 60 -38
rect 54 -48 60 -42
<< pdiffusion >>
rect 4 0 10 2
rect 4 -4 5 0
rect 9 -4 10 0
rect 4 -18 10 -4
rect 12 0 27 2
rect 12 -4 13 0
rect 17 -4 27 0
rect 12 -18 27 -4
rect 29 0 36 2
rect 29 -4 30 0
rect 34 -4 36 0
rect 29 -18 36 -4
rect 46 -3 52 2
rect 46 -7 47 -3
rect 51 -7 52 -3
rect 46 -18 52 -7
rect 54 -3 60 2
rect 54 -7 55 -3
rect 59 -7 60 -3
rect 54 -18 60 -7
<< metal1 >>
rect 4 12 70 13
rect 4 8 5 12
rect 9 8 30 12
rect 34 10 70 12
rect 34 8 47 10
rect 4 6 47 8
rect 51 6 70 10
rect 4 5 70 6
rect 5 0 9 5
rect 30 0 34 5
rect 47 -3 51 5
rect 13 -21 17 -4
rect 13 -23 39 -21
rect 13 -25 48 -23
rect 35 -27 48 -25
rect 35 -37 39 -27
rect 17 -41 22 -37
rect 34 -41 39 -37
rect 55 -38 59 -7
rect 5 -51 9 -41
rect 47 -51 51 -42
rect 5 -53 71 -51
rect 5 -54 47 -53
rect 9 -57 47 -54
rect 51 -57 71 -53
rect 9 -58 71 -57
rect 5 -61 71 -58
<< ntransistor >>
rect 10 -48 12 -36
rect 27 -48 29 -36
rect 52 -48 54 -30
<< ptransistor >>
rect 10 -18 12 2
rect 27 -18 29 2
rect 52 -18 54 2
<< polycontact >>
rect 6 -28 10 -24
rect 23 -32 27 -28
rect 48 -27 52 -23
<< ndcontact >>
rect 5 -41 9 -37
rect 13 -41 17 -37
rect 22 -41 26 -37
rect 30 -41 34 -37
rect 47 -42 51 -38
rect 55 -42 59 -38
<< pdcontact >>
rect 5 -4 9 0
rect 13 -4 17 0
rect 30 -4 34 0
rect 47 -7 51 -3
rect 55 -7 59 -3
<< psubstratepcontact >>
rect 5 -58 9 -54
rect 47 -57 51 -53
<< nsubstratencontact >>
rect 5 8 9 12
rect 30 8 34 12
rect 47 6 51 10
<< labels >>
rlabel metal1 57 -25 57 -25 1 out
rlabel metal1 63 9 63 9 5 Vdd
rlabel metal1 64 -56 64 -56 1 Vss
rlabel polycontact 26 -30 26 -30 1 b
rlabel polycontact 8 -26 8 -26 3 a
<< end >>
