* SPICE3 file created from nand2.ext - technology: scmos

.option scale=1u

M1000 out a Vdd Vdd pfet w=20 l=2
+  ad=300 pd=70 as=120 ps=52
M1001 a_12_13# a Vss Gnd nfet w=12 l=2
+  ad=144 pd=72 as=72 ps=36
M1002 out b a_12_13# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1003 a_29_43# b out Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 Vss Gnd 13.44fF
C1 out Gnd 4.61fF
C2 b Gnd 6.27fF
C3 a Gnd 6.27fF
